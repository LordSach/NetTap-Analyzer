// ************************************************************************************************************************
//
// PROJECT      :   NetTap-Analyzer
// PRODUCT      :   NetTap-DMA
// FILE         :   mm2s_top.sv
// AUTHOR       :   Sachith Rathnayake
// DESCRIPTION  :   mm2s_top module of DMA core
//
// ************************************************************************************************************************
//
// REVISIONS:
//
//  Date           Developer               Description
//  -----------    --------------------    -----------
//  19-Nov-2025    Sachith Rathnayake      Design
//
//
//*************************************************************************************************************************

`timescale 1ns/1ps

module mm2s_top (
    clk,
    rst_n,

    // AXI-MM Read
    m_axi_araddr,
    m_axi_arlen,
    m_axi_arvalid,
    m_axi_arready,
    m_axi_rdata,
    m_axi_rvalid,
    m_axi_rready,
    m_axi_rlast,

    // AXI-Stream Out
    m_axis_tdata,
    m_axis_tkeep,
    m_axis_tvalid,
    m_axis_tready,
    m_axis_tlast
);

    //---------------------------------------------------------------------------------------------------------------------
    // Global constant headers
    //---------------------------------------------------------------------------------------------------------------------
    
    
    
    //---------------------------------------------------------------------------------------------------------------------
    // parameter definitions
    //---------------------------------------------------------------------------------------------------------------------
    
    
    
    //---------------------------------------------------------------------------------------------------------------------
    // localparam definitions
    //---------------------------------------------------------------------------------------------------------------------
    
    
    
    //---------------------------------------------------------------------------------------------------------------------
    // type definitions
    //---------------------------------------------------------------------------------------------------------------------
    
    
    
    //---------------------------------------------------------------------------------------------------------------------
    // I/O signals
    //---------------------------------------------------------------------------------------------------------------------
    // Clock and negative reset
    input   logic           clk;
    input   logic           rst_n;

    // AXI-MM Read
    output  logic [31:0]    m_axi_araddr;
    output  logic [7:0]     m_axi_arlen;
    output  logic           m_axi_arvalid;
    input   logic           m_axi_arready;
    input   logic [31:0]    m_axi_rdata;
    input   logic           m_axi_rvalid;
    output  logic           m_axi_rready;
    input   logic           m_axi_rlast;

    // AXI-Stream Out
    output  logic [31:0]    m_axis_tdata;
    output  logic [3:0]     m_axis_tkeep;
    output  logic           m_axis_tvalid;
    input   logic           m_axis_tready;
    output  logic           m_axis_tlast;
    
    
    //---------------------------------------------------------------------------------------------------------------------
    // Internal signals
    //---------------------------------------------------------------------------------------------------------------------
    
    
    
    //---------------------------------------------------------------------------------------------------------------------
    // Implementation
    //---------------------------------------------------------------------------------------------------------------------
    
    
    
endmodule